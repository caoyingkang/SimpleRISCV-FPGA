module alu32(input      [31:0] srca,
             input      [31:0] srcb,
             input      [3:0]  alucontrol,
             input      [4:0]  shamt,
             output reg [31:0] aluresult,
             output            zero);

  wire [31:0] addresult;
  wire        sub, slt;

  lookahead_adder32 src_add(srca, srcb, sub, addresult);

  assign sub = alucontrol[3] | (~alucontrol[2] & alucontrol[1]);
  assign slt = (srca[31] & ~srcb[31]) |
               (srca[31] & srcb[31] & addresult[31]) |
               (~srca[31] & ~srcb[31] & addresult[31]);
  assign zero = (addresult == 32'b0);

  always @( * )
  begin
    case(alucontrol[2:0])
      3'b000:  aluresult = addresult; // ADD/SUB/ADDI.
      3'b001:  aluresult = srca << shamt; // SLLI. unimplemented:SLL.
      3'b010:  aluresult = slt; // SLT/SLTI
      3'b011:  aluresult = {32{1'bx}}; // unimplemented:SLTU/SLTIU.
      3'b100:  aluresult = srca ^ srcb; // XOR/XORI
      3'b101:  aluresult = {{1'b0}, srca[31:1]}; // SRLI (only shift by 1 in this lab). unimplemented: SRL/SRA/SRAI
      3'b110:  aluresult = srca | srcb; // OR/ORI
      3'b111:  aluresult = srca & srcb; // AND/ANDI
      default: aluresult = {(32){1'bx}};
    endcase
  end
endmodule

module lookahead_adder32(input  [31:0] srca,
                         input  [31:0] srcb,
                         input         sub,
                         output [31:0] addresult);

  wire [31:0] g, p, c, srcbneg, srcbadd;

  mux2 #(32) add_or_sub(srcb, srcbneg, sub, srcbadd);

  assign srcbneg = ~srcb;
  assign g = srca & srcbadd;
  assign p = srca ^ srcbadd;
  assign addresult = p ^ c;

  assign c[0] = sub;
  assign c[1] = g[0]
              | (p[0] & sub);
  assign c[2] = g[1]
              | (p[1] & g[0]) 
              | (p[1] & p[0] & sub);
  assign c[3] = g[2]
              | (p[2] & g[1]) 
              | (p[2] & p[1] & g[0]) 
              | (p[2] & p[1] & p[0] & sub);
  assign c[4] = g[3]
              | (p[3] & g[2]) 
              | (p[3] & p[2] & g[1]) 
              | (p[3] & p[2] & p[1] & g[0]) 
              | (p[3] & p[2] & p[1] & p[0] & sub);
  assign c[5] = g[4] 
              | (p[4] & g[3]) 
              | (p[4] & p[3] & g[2]) 
              | (p[4] & p[3] & p[2] & g[1]) 
              | (p[4] & p[3] & p[2] & p[1] & g[0]) 
              | (p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[6] = g[5] 
              | (p[5] & g[4]) 
              | (p[5] & p[4] & g[3]) 
              | (p[5] & p[4] & p[3] & g[2])
              | (p[5] & p[4] & p[3] & p[2] & g[1]) 
              | (p[5] & p[4] & p[3] & p[2] & p[1] & g[0]) 
              | (p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[7] = g[6]
              | (p[6] & g[5]) 
              | (p[6] & p[5] & g[4]) 
              | (p[6] & p[5] & p[4] & g[3]) 
              | (p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) 
              | (p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0]) 
              | (p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[8] = g[7]
              | (p[7] & g[6])
              | (p[7] & p[6] & g[5]) 
              | (p[7] & p[6] & p[5] & g[4]) 
              | (p[7] & p[6] & p[5] & p[4] & g[3]) 
              | (p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) 
              | (p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0]) 
              | (p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[9] = g[8]
              | (p[8] & g[7])
              | (p[8] & p[7] & g[6])
              | (p[8] & p[7] & p[6] & g[5]) 
              | (p[8] & p[7] & p[6] & p[5] & g[4]) 
              | (p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) 
              | (p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) 
              | (p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0]) 
              | (p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[10] = g[9]
              | (p[9] & g[8])
              | (p[9] & p[8] & g[7])
              | (p[9] & p[8] & p[7] & g[6])
              | (p[9] & p[8] & p[7] & p[6] & g[5]) 
              | (p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) 
              | (p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) 
              | (p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) 
              | (p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0]) 
              | (p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[11] = g[10]
              | (p[10] & g[9])
              | (p[10] & p[9] & g[8])
              | (p[10] & p[9] & p[8] & g[7])
              | (p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) 
              | (p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) 
              | (p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) 
              | (p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) 
              | (p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0]) 
              | (p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[12] = g[11]
              | (p[11] & g[10])
              | (p[11] & p[10] & g[9])
              | (p[11] & p[10] & p[9] & g[8])
              | (p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[13] = g[12]
              | (p[12] & g[11])
              | (p[12] & p[11] & g[10])
              | (p[12] & p[11] & p[10] & g[9])
              | (p[12] & p[11] & p[10] & p[9] & g[8])
              | (p[12] & p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[14] = g[13]
              | (p[13] & g[12])
              | (p[13] & p[12] & g[11])
              | (p[13] & p[12] & p[11] & g[10])
              | (p[13] & p[12] & p[11] & p[10] & g[9])
              | (p[13] & p[12] & p[11] & p[10] & p[9] & g[8])
              | (p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[15] = g[14]
              | (p[14] & g[13])
              | (p[14] & p[13] & g[12])
              | (p[14] & p[13] & p[12] & g[11])
              | (p[14] & p[13] & p[12] & p[11] & g[10])
              | (p[14] & p[13] & p[12] & p[11] & p[10] & g[9])
              | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8])
              | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[16] = g[15]
              | (p[15] & g[14])
              | (p[15] & p[14] & g[13])
              | (p[15] & p[14] & p[13] & g[12])
              | (p[15] & p[14] & p[13] & p[12] & g[11])
              | (p[15] & p[14] & p[13] & p[12] & p[11] & g[10])
              | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9])
              | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8])
              | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[17] = g[16]
              | (p[16] & g[15])
              | (p[16] & p[15] & g[14])
              | (p[16] & p[15] & p[14] & g[13])
              | (p[16] & p[15] & p[14] & p[13] & g[12])
              | (p[16] & p[15] & p[14] & p[13] & p[12] & g[11])
              | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10])
              | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9])
              | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8])
              | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[18] = g[17]
              | (p[17] & g[16])
              | (p[17] & p[16] & g[15])
              | (p[17] & p[16] & p[15] & g[14])
              | (p[17] & p[16] & p[15] & p[14] & g[13])
              | (p[17] & p[16] & p[15] & p[14] & p[13] & g[12])
              | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11])
              | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10])
              | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9])
              | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8])
              | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[19] = g[18]
              | (p[18] & g[17])
              | (p[18] & p[17] & g[16])
              | (p[18] & p[17] & p[16] & g[15])
              | (p[18] & p[17] & p[16] & p[15] & g[14])
              | (p[18] & p[17] & p[16] & p[15] & p[14] & g[13])
              | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12])
              | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11])
              | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10])
              | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9])
              | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8])
              | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[20] = g[19]
              | (p[19] & g[18])
              | (p[19] & p[18] & g[17])
              | (p[19] & p[18] & p[17] & g[16])
              | (p[19] & p[18] & p[17] & p[16] & g[15])
              | (p[19] & p[18] & p[17] & p[16] & p[15] & g[14])
              | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13])
              | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12])
              | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11])
              | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10])
              | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9])
              | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8])
              | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[21] = g[20]
              | (p[20] & g[19])
              | (p[20] & p[19] & g[18])
              | (p[20] & p[19] & p[18] & g[17])
              | (p[20] & p[19] & p[18] & p[17] & g[16])
              | (p[20] & p[19] & p[18] & p[17] & p[16] & g[15])
              | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14])
              | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13])
              | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12])
              | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11])
              | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10])
              | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9])
              | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8])
              | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[22] = g[21]
              | (p[21] & g[20])
              | (p[21] & p[20] & g[19])
              | (p[21] & p[20] & p[19] & g[18])
              | (p[21] & p[20] & p[19] & p[18] & g[17])
              | (p[21] & p[20] & p[19] & p[18] & p[17] & g[16])
              | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15])
              | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14])
              | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13])
              | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12])
              | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11])
              | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10])
              | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9])
              | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8])
              | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[23] = g[22]
              | (p[22] & g[21])
              | (p[22] & p[21] & g[20])
              | (p[22] & p[21] & p[20] & g[19])
              | (p[22] & p[21] & p[20] & p[19] & g[18])
              | (p[22] & p[21] & p[20] & p[19] & p[18] & g[17])
              | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & g[16])
              | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15])
              | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14])
              | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13])
              | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12])
              | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11])
              | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10])
              | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9])
              | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8])
              | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[24] = g[23]
              | (p[23] & g[22])
              | (p[23] & p[22] & g[21])
              | (p[23] & p[22] & p[21] & g[20])
              | (p[23] & p[22] & p[21] & p[20] & g[19])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & g[18])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & g[17])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & g[16])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[25] = g[24]
              | (p[24] & g[23])
              | (p[24] & p[23] & g[22])
              | (p[24] & p[23] & p[22] & g[21])
              | (p[24] & p[23] & p[22] & p[21] & g[20])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & g[19])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & g[18])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & g[17])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & g[16])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[26] = g[25]
              | (p[25] & g[24])
              | (p[25] & p[24] & g[23])
              | (p[25] & p[24] & p[23] & g[22])
              | (p[25] & p[24] & p[23] & p[22] & g[21])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & g[20])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & g[19])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & g[18])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & g[17])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & g[16])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[27] = g[26]
              | (p[26] & g[25])
              | (p[26] & p[25] & g[24])
              | (p[26] & p[25] & p[24] & g[23])
              | (p[26] & p[25] & p[24] & p[23] & g[22])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & g[21])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & g[20])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & g[19])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & g[18])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & g[17])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & g[16])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[28] = g[27]
              | (p[27] & g[26])
              | (p[27] & p[26] & g[25])
              | (p[27] & p[26] & p[25] & g[24])
              | (p[27] & p[26] & p[25] & p[24] & g[23])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & g[22])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & g[21])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & g[20])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & g[19])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & g[18])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & g[17])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & g[16])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[29] = g[28]
              | (p[28] & g[27])
              | (p[28] & p[27] & g[26])
              | (p[28] & p[27] & p[26] & g[25])
              | (p[28] & p[27] & p[26] & p[25] & g[24])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & g[23])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & g[22])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & g[21])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & g[20])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & g[19])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & g[18])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & g[17])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & g[16])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[30] = g[29]
              | (p[29] & g[28])
              | (p[29] & p[28] & g[27])
              | (p[29] & p[28] & p[27] & g[26])
              | (p[29] & p[28] & p[27] & p[26] & g[25])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & g[24])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & g[23])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & g[22])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & g[21])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & g[20])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & g[19])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & g[18])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & g[17])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & g[16])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
  assign c[31] = g[30]
              | (p[30] & g[29])
              | (p[30] & p[29] & g[28])
              | (p[30] & p[29] & p[28] & g[27])
              | (p[30] & p[29] & p[28] & p[27] & g[26])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & g[25])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & g[24])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & g[23])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & g[22])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & g[21])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & g[20])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & g[19])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & g[18])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & g[17])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & g[16])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])
              | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & p[0] & sub);
endmodule